class baseClass;
	int data;
	function new();
		data=32'hc0de_c0de;
	endfuction
endclass
